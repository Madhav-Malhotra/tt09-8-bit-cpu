/*
 * Copyright (c) 2024 WAT.ai Chip Team
 * SPDX-License-Identifier: Apache-2.0
 * Implements register A
 */

`include "../common/bus_transceiver.v"

module regA_top (
    input wire clk,
    input wire [7:0] bus,
    input wire clr,
    input wire ai_n,
    input wire ao_n,
    output wire [7:0] A
);

    

endmodule